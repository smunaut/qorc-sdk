/*
 * s3_inc8.v
 *
 * vim: ts=4 sw=4
 *
 * Combinatorial 8-bit incrementer implemented in 5 LCs with 2 layers
 * of logic.
 *
 * Copyright (C) 2020 Sylvain Munaut
 * All rights reserved.
 *
 * LGPL v3+, see LICENSE.lgpl3
 *
 * This program is free software; you can redistribute it and/or
 * modify it under the terms of the GNU Lesser General Public
 * License as published by the Free Software Foundation; either
 * version 3 of the License, or (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
 * Lesser General Public License for more details.
 *
 * You should have received a copy of the GNU Lesser General Public License
 * along with this program; if not, write to the Free Software Foundation,
 * Inc., 51 Franklin Street, Fifth Floor, Boston, MA 02110-1301, USA.
 */

`default_nettype none

module s3_inc8 (
	input  wire [7:0] a,
	output wire [7:0] x
);

	wire carry;	// Carry generated by [3:0]
	wire a4_n;	// !a[4]
	wire int6;
	wire int7;

	// Cell 0
	//  - bit [0] using FMUX   (FZ out)
	//  - bit [1] using Bottom (CZ out)
	//  - bit [2] using Top    (TZ out)

	logic_cell_macro cell_0_I (
		.BA1  (1'b0),	// 00
		.BA2  (1'b1),	// 10
		.BAB  (a[0]),
		.BAS1 (1'b0),
		.BAS2 (1'b0),
		.BB1  (1'b1),	// 01
		.BB2  (1'b0),	// 11
		.BBS1 (1'b0),
		.BBS2 (1'b0),
		.BSL  (a[1]),
		.F1   (1'b1),
		.F2   (1'b0),
		.FS   (a[0]),
		.QCK  (1'b0),
		.QCKS (1'b0),
		.QDI  (1'b0),
		.QDS  (1'b0),
		.QEN  (1'b0),
		.QRT  (1'b0),
		.QST  (1'b0),
		.TA1  (a[2]),
		.TA2  (a[2]),
		.TAB  (a[0]),
		.TAS1 (1'b0),
		.TAS2 (1'b0),
		.TB1  (a[2]),
		.TB2  (a[2]),
		.TBS  (1'b1),
		.TBS1 (1'b0),
		.TBS2 (1'b1),
		.TSL  (a[1]),
		.CZ   (x[1]),
		.FZ   (x[0]),
		.QZ   (),
		.TZ   (x[2])
	);


	// Cell 1
	//  - pre bit [4] invert using FMUX (FZ out)
	//  - bit [3] using LUT4 (CZ out)

	logic_cell_macro cell_1_I (
		.BA1  (a[3]),
		.BA2  (a[3]),
		.BAB  (a[0]),
		.BAS1 (1'b0),
		.BAS2 (1'b0),
		.BB1  (a[3]),
		.BB2  (a[3]),
		.BBS1 (1'b0),
		.BBS2 (1'b1),
		.BSL  (a[1]),
		.F1   (1'b1),
		.F2   (1'b0),
		.FS   (a[4]),
		.QCK  (1'b0),
		.QCKS (1'b0),
		.QDI  (1'b0),
		.QDS  (1'b0),
		.QEN  (1'b0),
		.QRT  (1'b0),
		.QST  (1'b0),
		.TA1  (a[3]),
		.TA2  (1'b0),
		.TAB  (1'b0),
		.TAS1 (1'b0),
		.TAS2 (1'b0),
		.TB1  (1'b0),
		.TB2  (1'b0),
		.TBS  (a[2]),
		.TBS1 (1'b0),
		.TBS2 (1'b0),
		.TSL  (1'b0),
		.CZ   (x[3]),
		.FZ   (a4_n),
		.QZ   (),
		.TZ   ()
	);


	// Cell 2
	//  - bit [4] using FMUX (FZ out)
	//  - carry gen using LUT4 (CZ out)

	logic_cell_macro cell_2_I (
		.BA1  (1'b0),
		.BA2  (1'b0),
		.BAB  (a[0]),
		.BAS1 (1'b0),
		.BAS2 (1'b0),
		.BB1  (1'b0),
		.BB2  (a[3]),
		.BBS1 (1'b0),
		.BBS2 (1'b0),
		.BSL  (a[1]),
		.F1   (a[4]),
		.F2   (a4_n),
		.FS   (carry),
		.QCK  (1'b0),
		.QCKS (1'b0),
		.QDI  (1'b0),
		.QDS  (1'b0),
		.QEN  (1'b0),
		.QRT  (1'b0),
		.QST  (1'b0),
		.TA1  (1'b0),
		.TA2  (1'b0),
		.TAB  (1'b0),
		.TAS1 (1'b0),
		.TAS2 (1'b0),
		.TB1  (1'b0),
		.TB2  (1'b0),
		.TBS  (a[2]),
		.TBS1 (1'b0),
		.TBS2 (1'b0),
		.TSL  (1'b0),
		.CZ   (carry),
		.FZ   (x[4]),
		.QZ   (),
		.TZ   ()
	);

	// Cell 3
	//  - bit[5] using Top (TZ out)
	//  - bit[6] using Bottom + FMUX (FZ out)

	logic_cell_macro cell_3_I (
		.BA1  (a[6]),
		.BA2  (a[6]),
		.BAB  (a[4]),
		.BAS1 (1'b0),
		.BAS2 (1'b0),
		.BB1  (a[6]),
		.BB2  (a[6]),
		.BBS1 (1'b0),
		.BBS2 (1'b1),
		.BSL  (a[5]),
		.F1   (a[6]),
		.F2   (int6),
		.FS   (carry),
		.QCK  (1'b0),
		.QCKS (1'b0),
		.QDI  (1'b0),
		.QDS  (1'b0),
		.QEN  (1'b0),
		.QRT  (1'b0),
		.QST  (1'b0),
		.TA1  (1'b0),
		.TA2  (1'b1),
		.TAB  (carry),
		.TAS1 (1'b0),
		.TAS2 (1'b0),
		.TB1  (a[4]),
		.TB2  (a[4]),
		.TBS  (1'b1),
		.TBS1 (1'b0),
		.TBS2 (1'b1),
		.TSL  (a[5]),
		.CZ   (int6),
		.FZ   (x[6]),
		.QZ   (),
		.TZ   (x[5])
	);


	// Cell 4
	//  - bit[7] using LUT4 + FMUX (FZ out)

	logic_cell_macro cell_4_I (
		.BA1  (a[7]),
		.BA2  (a[7]),
		.BAB  (a[4]),
		.BAS1 (1'b0),
		.BAS2 (1'b0),
		.BB1  (a[7]),
		.BB2  (a[7]),
		.BBS1 (1'b0),
		.BBS2 (1'b1),
		.BSL  (a[5]),
		.F1   (a[7]),
		.F2   (int7),
		.FS   (carry),
		.QCK  (1'b0),
		.QCKS (1'b0),
		.QDI  (1'b0),
		.QDS  (1'b0),
		.QEN  (1'b0),
		.QRT  (1'b0),
		.QST  (1'b0),
		.TA1  (a[7]),
		.TA2  (1'b0),
		.TAB  (1'b0),
		.TAS1 (1'b0),
		.TAS2 (1'b0),
		.TB1  (1'b0),
		.TB2  (1'b0),
		.TBS  (a[6]),
		.TBS1 (1'b0),
		.TBS2 (1'b0),
		.TSL  (1'b0),
		.CZ   (int7),
		.FZ   (x[7]),
		.QZ   (),
		.TZ   ()
	);

endmodule // s3_inc8
